module ShiftRight(
  input  [4:0] io_in,
  output [4:0] io_out
);
  assign io_out = {{3'd0}, io_in[4:3]}; // @[ArithmeticLogical.scala 103:21]
endmodule
module ShiftRight_1(
  input  [12:0] io_in,
  output [12:0] io_out
);
  assign io_out = {{4'd0}, io_in[12:4]}; // @[ArithmeticLogical.scala 103:21]
endmodule
module RandomHardware_1_1(
  input  [12:0] io_in,
  output [12:0] io_out
);
  wire [12:0] ShiftRight_000_io_in; // @[RandomHardware_1_1.scala 14:34]
  wire [12:0] ShiftRight_000_io_out; // @[RandomHardware_1_1.scala 14:34]
  ShiftRight_1 ShiftRight_000 ( // @[RandomHardware_1_1.scala 14:34]
    .io_in(ShiftRight_000_io_in),
    .io_out(ShiftRight_000_io_out)
  );
  assign io_out = ShiftRight_000_io_out; // @[RandomHardware_1_1.scala 17:10]
  assign ShiftRight_000_io_in = io_in; // @[RandomHardware_1_1.scala 16:25]
endmodule
module Accum(
  input        clock,
  input  [7:0] io_in,
  output [7:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] sum; // @[ArithmeticLogical.scala 82:18]
  assign io_out = sum; // @[ArithmeticLogical.scala 84:12]
  always @(posedge clock) begin
    sum <= sum + io_in; // @[ArithmeticLogical.scala 83:16]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sum = _RAND_0[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ReduceXorMux(
  input  [19:0] io_in,
  output [7:0]  io_out
);
  wire [7:0] IN1 = io_in[19:12]; // @[Muxes.scala 122:27]
  wire [7:0] IN2 = io_in[11:4]; // @[Muxes.scala 123:27]
  wire [3:0] SEL = io_in[3:0]; // @[Muxes.scala 124:27]
  assign io_out = ^SEL ? IN1 : IN2; // @[Muxes.scala 126:18]
endmodule
module RandomHardware_2_0(
  input         clock,
  input  [19:0] io_in,
  output [7:0]  io_out
);
  wire  Accum_000_clock; // @[RandomHardware_2_0.scala 15:34]
  wire [7:0] Accum_000_io_in; // @[RandomHardware_2_0.scala 15:34]
  wire [7:0] Accum_000_io_out; // @[RandomHardware_2_0.scala 15:34]
  wire [19:0] ReduceXorMux_001_io_in; // @[RandomHardware_2_0.scala 16:34]
  wire [7:0] ReduceXorMux_001_io_out; // @[RandomHardware_2_0.scala 16:34]
  Accum Accum_000 ( // @[RandomHardware_2_0.scala 15:34]
    .clock(Accum_000_clock),
    .io_in(Accum_000_io_in),
    .io_out(Accum_000_io_out)
  );
  ReduceXorMux ReduceXorMux_001 ( // @[RandomHardware_2_0.scala 16:34]
    .io_in(ReduceXorMux_001_io_in),
    .io_out(ReduceXorMux_001_io_out)
  );
  assign io_out = Accum_000_io_out; // @[RandomHardware_2_0.scala 19:10]
  assign Accum_000_clock = clock;
  assign Accum_000_io_in = ReduceXorMux_001_io_out; // @[RandomHardware_2_0.scala 13:24 RandomHardware_2_0.scala 21:18]
  assign ReduceXorMux_001_io_in = io_in; // @[RandomHardware_2_0.scala 18:33]
endmodule
module RegE(
  input         clock,
  input  [19:0] io_in,
  output [18:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [18:0] data = io_in[19:1]; // @[Memory.scala 20:21]
  wire  en = io_in[0]; // @[Memory.scala 21:19]
  reg [17:0] reg_; // @[Memory.scala 22:18]
  wire [18:0] _GEN_0 = en ? data : {{1'd0}, reg_}; // @[Memory.scala 23:14 Memory.scala 23:20 Memory.scala 22:18]
  assign io_out = {{1'd0}, reg_}; // @[Memory.scala 24:12]
  always @(posedge clock) begin
    reg_ <= _GEN_0[17:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_ = _RAND_0[17:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RandomHardware_2_1(
  input         clock,
  input  [19:0] io_in,
  output [18:0] io_out
);
  wire  RegE_000_clock; // @[RandomHardware_2_1.scala 14:26]
  wire [19:0] RegE_000_io_in; // @[RandomHardware_2_1.scala 14:26]
  wire [18:0] RegE_000_io_out; // @[RandomHardware_2_1.scala 14:26]
  RegE RegE_000 ( // @[RandomHardware_2_1.scala 14:26]
    .clock(RegE_000_clock),
    .io_in(RegE_000_io_in),
    .io_out(RegE_000_io_out)
  );
  assign io_out = RegE_000_io_out; // @[RandomHardware_2_1.scala 17:10]
  assign RegE_000_clock = clock;
  assign RegE_000_io_in = io_in; // @[RandomHardware_2_1.scala 16:25]
endmodule
module RandomHardware_1_3(
  input         clock,
  input  [15:0] io_in,
  output [17:0] io_out
);
  wire  RandomHardware_000_clock; // @[RandomHardware_1_3.scala 15:42]
  wire [19:0] RandomHardware_000_io_in; // @[RandomHardware_1_3.scala 15:42]
  wire [7:0] RandomHardware_000_io_out; // @[RandomHardware_1_3.scala 15:42]
  wire  RandomHardware_001_clock; // @[RandomHardware_1_3.scala 16:42]
  wire [19:0] RandomHardware_001_io_in; // @[RandomHardware_1_3.scala 16:42]
  wire [18:0] RandomHardware_001_io_out; // @[RandomHardware_1_3.scala 16:42]
  wire [14:0] wire_000 = {{7'd0}, RandomHardware_000_io_out}; // @[RandomHardware_1_3.scala 13:24 RandomHardware_1_3.scala 21:18]
  RandomHardware_2_0 RandomHardware_000 ( // @[RandomHardware_1_3.scala 15:42]
    .clock(RandomHardware_000_clock),
    .io_in(RandomHardware_000_io_in),
    .io_out(RandomHardware_000_io_out)
  );
  RandomHardware_2_1 RandomHardware_001 ( // @[RandomHardware_1_3.scala 16:42]
    .clock(RandomHardware_001_clock),
    .io_in(RandomHardware_001_io_in),
    .io_out(RandomHardware_001_io_out)
  );
  assign io_out = RandomHardware_001_io_out[17:0]; // @[RandomHardware_1_3.scala 19:10]
  assign RandomHardware_000_clock = clock;
  assign RandomHardware_000_io_in = {{4'd0}, io_in}; // @[RandomHardware_1_3.scala 18:33]
  assign RandomHardware_001_clock = clock;
  assign RandomHardware_001_io_in = {{5'd0}, wire_000}; // @[RandomHardware_1_3.scala 13:24 RandomHardware_1_3.scala 21:18]
endmodule
module SignExtendDouble(
  input  [14:0] io_in,
  output [29:0] io_out
);
  wire [14:0] io_out_hi = io_in[14] ? 15'h7fff : 15'h0; // @[Bitwise.scala 72:12]
  assign io_out = {io_out_hi,io_in}; // @[Cat.scala 30:58]
endmodule
module Reg(
  input         clock,
  input  [36:0] io_in,
  output [36:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [36:0] io_out_REG; // @[Memory.scala 12:22]
  assign io_out = io_out_REG; // @[Memory.scala 12:12]
  always @(posedge clock) begin
    io_out_REG <= io_in; // @[Memory.scala 12:22]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  io_out_REG = _RAND_0[36:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RandomHardware_1_4(
  input         clock,
  input  [36:0] io_in,
  output [29:0] io_out
);
  wire [14:0] SignExtendDouble_000_io_in; // @[RandomHardware_1_4.scala 16:42]
  wire [29:0] SignExtendDouble_000_io_out; // @[RandomHardware_1_4.scala 16:42]
  wire  RandomHardware_001_clock; // @[RandomHardware_1_4.scala 17:42]
  wire [19:0] RandomHardware_001_io_in; // @[RandomHardware_1_4.scala 17:42]
  wire [18:0] RandomHardware_001_io_out; // @[RandomHardware_1_4.scala 17:42]
  wire  Reg_002_clock; // @[RandomHardware_1_4.scala 18:26]
  wire [36:0] Reg_002_io_in; // @[RandomHardware_1_4.scala 18:26]
  wire [36:0] Reg_002_io_out; // @[RandomHardware_1_4.scala 18:26]
  wire [36:0] wire_001 = Reg_002_io_out; // @[RandomHardware_1_4.scala 14:24 RandomHardware_1_4.scala 25:18]
  SignExtendDouble SignExtendDouble_000 ( // @[RandomHardware_1_4.scala 16:42]
    .io_in(SignExtendDouble_000_io_in),
    .io_out(SignExtendDouble_000_io_out)
  );
  RandomHardware_2_1 RandomHardware_001 ( // @[RandomHardware_1_4.scala 17:42]
    .clock(RandomHardware_001_clock),
    .io_in(RandomHardware_001_io_in),
    .io_out(RandomHardware_001_io_out)
  );
  Reg Reg_002 ( // @[RandomHardware_1_4.scala 18:26]
    .clock(Reg_002_clock),
    .io_in(Reg_002_io_in),
    .io_out(Reg_002_io_out)
  );
  assign io_out = SignExtendDouble_000_io_out; // @[RandomHardware_1_4.scala 21:10]
  assign SignExtendDouble_000_io_in = RandomHardware_001_io_out[14:0]; // @[RandomHardware_1_4.scala 13:24 RandomHardware_1_4.scala 24:18]
  assign RandomHardware_001_clock = clock;
  assign RandomHardware_001_io_in = wire_001[19:0]; // @[RandomHardware_1_4.scala 23:33]
  assign Reg_002_clock = clock;
  assign Reg_002_io_in = io_in; // @[RandomHardware_1_4.scala 20:25]
endmodule
module ShiftRegister(
  input        clock,
  input  [4:0] io_in,
  output [4:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] r0; // @[Memory.scala 78:19]
  reg [4:0] r1; // @[Memory.scala 79:19]
  reg [4:0] r2; // @[Memory.scala 80:19]
  reg [4:0] r3; // @[Memory.scala 81:19]
  assign io_out = r3; // @[Memory.scala 82:10]
  always @(posedge clock) begin
    r0 <= io_in; // @[Memory.scala 78:19]
    r1 <= r0; // @[Memory.scala 79:19]
    r2 <= r1; // @[Memory.scala 80:19]
    r3 <= r2; // @[Memory.scala 81:19]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r0 = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  r1 = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  r2 = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  r3 = _RAND_3[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Reg_1(
  input        clock,
  input  [7:0] io_in,
  output [7:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] io_out_REG; // @[Memory.scala 12:22]
  assign io_out = io_out_REG; // @[Memory.scala 12:12]
  always @(posedge clock) begin
    io_out_REG <= io_in; // @[Memory.scala 12:22]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  io_out_REG = _RAND_0[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SignExtendDouble_1(
  input  [9:0]  io_in,
  output [19:0] io_out
);
  wire [9:0] io_out_hi = io_in[9] ? 10'h3ff : 10'h0; // @[Bitwise.scala 72:12]
  assign io_out = {io_out_hi,io_in}; // @[Cat.scala 30:58]
endmodule
module Mux2(
  input  [20:0] io_in,
  output [9:0]  io_out
);
  wire  sel = io_in[20]; // @[Muxes.scala 16:18]
  wire [9:0] in1 = io_in[19:10]; // @[Muxes.scala 17:18]
  wire [9:0] in0 = io_in[9:0]; // @[Muxes.scala 18:18]
  assign io_out = sel ? in1 : in0; // @[Muxes.scala 19:15 Muxes.scala 19:24 Muxes.scala 20:24]
endmodule
module RandomHardware_2_2(
  input  [20:0] io_in,
  output [9:0]  io_out
);
  wire [20:0] Mux2_000_io_in; // @[RandomHardware_2_2.scala 14:26]
  wire [9:0] Mux2_000_io_out; // @[RandomHardware_2_2.scala 14:26]
  Mux2 Mux2_000 ( // @[RandomHardware_2_2.scala 14:26]
    .io_in(Mux2_000_io_in),
    .io_out(Mux2_000_io_out)
  );
  assign io_out = Mux2_000_io_out; // @[RandomHardware_2_2.scala 17:10]
  assign Mux2_000_io_in = io_in; // @[RandomHardware_2_2.scala 16:25]
endmodule
module ShiftLeft(
  input  [18:0] io_in,
  output [22:0] io_out
);
  assign io_out = {io_in, 4'h0}; // @[ArithmeticLogical.scala 94:21]
endmodule
module RandomHardware_1_7(
  input         clock,
  input  [20:0] io_in,
  output [22:0] io_out
);
  wire [9:0] SignExtendDouble_000_io_in; // @[RandomHardware_1_7.scala 17:42]
  wire [19:0] SignExtendDouble_000_io_out; // @[RandomHardware_1_7.scala 17:42]
  wire  RandomHardware_001_clock; // @[RandomHardware_1_7.scala 18:42]
  wire [19:0] RandomHardware_001_io_in; // @[RandomHardware_1_7.scala 18:42]
  wire [18:0] RandomHardware_001_io_out; // @[RandomHardware_1_7.scala 18:42]
  wire [20:0] RandomHardware_002_io_in; // @[RandomHardware_1_7.scala 19:42]
  wire [9:0] RandomHardware_002_io_out; // @[RandomHardware_1_7.scala 19:42]
  wire [18:0] ShiftLeft_003_io_in; // @[RandomHardware_1_7.scala 20:34]
  wire [22:0] ShiftLeft_003_io_out; // @[RandomHardware_1_7.scala 20:34]
  SignExtendDouble_1 SignExtendDouble_000 ( // @[RandomHardware_1_7.scala 17:42]
    .io_in(SignExtendDouble_000_io_in),
    .io_out(SignExtendDouble_000_io_out)
  );
  RandomHardware_2_1 RandomHardware_001 ( // @[RandomHardware_1_7.scala 18:42]
    .clock(RandomHardware_001_clock),
    .io_in(RandomHardware_001_io_in),
    .io_out(RandomHardware_001_io_out)
  );
  RandomHardware_2_2 RandomHardware_002 ( // @[RandomHardware_1_7.scala 19:42]
    .io_in(RandomHardware_002_io_in),
    .io_out(RandomHardware_002_io_out)
  );
  ShiftLeft ShiftLeft_003 ( // @[RandomHardware_1_7.scala 20:34]
    .io_in(ShiftLeft_003_io_in),
    .io_out(ShiftLeft_003_io_out)
  );
  assign io_out = ShiftLeft_003_io_out; // @[RandomHardware_1_7.scala 23:10]
  assign SignExtendDouble_000_io_in = RandomHardware_002_io_out; // @[RandomHardware_1_7.scala 13:24 RandomHardware_1_7.scala 29:18]
  assign RandomHardware_001_clock = clock;
  assign RandomHardware_001_io_in = SignExtendDouble_000_io_out; // @[RandomHardware_1_7.scala 14:24 RandomHardware_1_7.scala 26:18]
  assign RandomHardware_002_io_in = io_in; // @[RandomHardware_1_7.scala 22:33]
  assign ShiftLeft_003_io_in = RandomHardware_001_io_out; // @[RandomHardware_1_7.scala 15:24 RandomHardware_1_7.scala 28:18]
endmodule
module CompareMux(
  input  [15:0] io_in,
  output [4:0]  io_out
);
  wire [7:0] IN1 = io_in[15:8]; // @[Muxes.scala 134:27]
  wire [4:0] IN2 = io_in[10:6]; // @[Muxes.scala 135:27]
  wire [2:0] SEL1 = io_in[5:3]; // @[Muxes.scala 136:27]
  wire [2:0] SEL2 = io_in[2:0]; // @[Muxes.scala 137:27]
  wire [7:0] _io_out_T_1 = SEL1 >= SEL2 ? IN1 : {{3'd0}, IN2}; // @[Muxes.scala 139:18]
  assign io_out = _io_out_T_1[4:0]; // @[Muxes.scala 139:12]
endmodule
module RandomHardware_1_8(
  input  [15:0] io_in,
  output [4:0]  io_out
);
  wire [15:0] CompareMux_000_io_in; // @[RandomHardware_1_8.scala 14:34]
  wire [4:0] CompareMux_000_io_out; // @[RandomHardware_1_8.scala 14:34]
  CompareMux CompareMux_000 ( // @[RandomHardware_1_8.scala 14:34]
    .io_in(CompareMux_000_io_in),
    .io_out(CompareMux_000_io_out)
  );
  assign io_out = CompareMux_000_io_out; // @[RandomHardware_1_8.scala 17:10]
  assign CompareMux_000_io_in = io_in; // @[RandomHardware_1_8.scala 16:25]
endmodule
module ShiftRegister_1(
  input        clock,
  input  [3:0] io_in,
  output [3:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] r0; // @[Memory.scala 78:19]
  reg [3:0] r1; // @[Memory.scala 79:19]
  reg [3:0] r2; // @[Memory.scala 80:19]
  reg [3:0] r3; // @[Memory.scala 81:19]
  assign io_out = r3; // @[Memory.scala 82:10]
  always @(posedge clock) begin
    r0 <= io_in; // @[Memory.scala 78:19]
    r1 <= r0; // @[Memory.scala 79:19]
    r2 <= r1; // @[Memory.scala 80:19]
    r3 <= r2; // @[Memory.scala 81:19]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r0 = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  r1 = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  r2 = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  r3 = _RAND_3[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Accum_2(
  input        clock,
  input  [5:0] io_in,
  output [5:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [5:0] sum; // @[ArithmeticLogical.scala 82:18]
  assign io_out = sum; // @[ArithmeticLogical.scala 84:12]
  always @(posedge clock) begin
    sum <= sum + io_in; // @[ArithmeticLogical.scala 83:16]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sum = _RAND_0[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RandomHardware_1_11(
  input         clock,
  input  [15:0] io_in,
  output [3:0]  io_out
);
  wire  RandomHardware_000_clock; // @[RandomHardware_1_11.scala 14:42]
  wire [19:0] RandomHardware_000_io_in; // @[RandomHardware_1_11.scala 14:42]
  wire [7:0] RandomHardware_000_io_out; // @[RandomHardware_1_11.scala 14:42]
  RandomHardware_2_0 RandomHardware_000 ( // @[RandomHardware_1_11.scala 14:42]
    .clock(RandomHardware_000_clock),
    .io_in(RandomHardware_000_io_in),
    .io_out(RandomHardware_000_io_out)
  );
  assign io_out = RandomHardware_000_io_out[3:0]; // @[RandomHardware_1_11.scala 17:10]
  assign RandomHardware_000_clock = clock;
  assign RandomHardware_000_io_in = {{4'd0}, io_in}; // @[RandomHardware_1_11.scala 16:33]
endmodule
module RandomHardware_1_12(
  input         clock,
  input  [11:0] io_in,
  output [11:0] io_out
);
  wire  RandomHardware_000_clock; // @[RandomHardware_1_12.scala 14:42]
  wire [19:0] RandomHardware_000_io_in; // @[RandomHardware_1_12.scala 14:42]
  wire [7:0] RandomHardware_000_io_out; // @[RandomHardware_1_12.scala 14:42]
  RandomHardware_2_0 RandomHardware_000 ( // @[RandomHardware_1_12.scala 14:42]
    .clock(RandomHardware_000_clock),
    .io_in(RandomHardware_000_io_in),
    .io_out(RandomHardware_000_io_out)
  );
  assign io_out = {{4'd0}, RandomHardware_000_io_out}; // @[RandomHardware_1_12.scala 17:10]
  assign RandomHardware_000_clock = clock;
  assign RandomHardware_000_io_in = {{8'd0}, io_in}; // @[RandomHardware_1_12.scala 16:33]
endmodule
module Mux2_1(
  input  [18:0] io_in,
  output [8:0]  io_out
);
  wire  sel = io_in[18]; // @[Muxes.scala 16:18]
  wire [8:0] in1 = io_in[17:9]; // @[Muxes.scala 17:18]
  wire [8:0] in0 = io_in[8:0]; // @[Muxes.scala 18:18]
  assign io_out = sel ? in1 : in0; // @[Muxes.scala 19:15 Muxes.scala 19:24 Muxes.scala 20:24]
endmodule
module RandomHardware_1_13(
  input  [18:0] io_in,
  output [8:0]  io_out
);
  wire [18:0] Mux2_000_io_in; // @[RandomHardware_1_13.scala 14:26]
  wire [8:0] Mux2_000_io_out; // @[RandomHardware_1_13.scala 14:26]
  Mux2_1 Mux2_000 ( // @[RandomHardware_1_13.scala 14:26]
    .io_in(Mux2_000_io_in),
    .io_out(Mux2_000_io_out)
  );
  assign io_out = Mux2_000_io_out; // @[RandomHardware_1_13.scala 17:10]
  assign Mux2_000_io_in = io_in; // @[RandomHardware_1_13.scala 16:25]
endmodule
module Mul(
  input  [5:0] io_in,
  output [5:0] io_out
);
  wire [2:0] in1 = io_in[5:3]; // @[ArithmeticLogical.scala 47:20]
  wire [2:0] in2 = io_in[2:0]; // @[ArithmeticLogical.scala 48:20]
  assign io_out = in1 * in2; // @[ArithmeticLogical.scala 49:19]
endmodule
module Reg_2(
  input        clock,
  input  [3:0] io_in,
  output [3:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] io_out_REG; // @[Memory.scala 12:22]
  assign io_out = io_out_REG; // @[Memory.scala 12:12]
  always @(posedge clock) begin
    io_out_REG <= io_in; // @[Memory.scala 12:22]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  io_out_REG = _RAND_0[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RegE_3(
  input         clock,
  input  [18:0] io_in,
  output [17:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [17:0] data = io_in[18:1]; // @[Memory.scala 20:21]
  wire  en = io_in[0]; // @[Memory.scala 21:19]
  reg [16:0] reg_; // @[Memory.scala 22:18]
  wire [17:0] _GEN_0 = en ? data : {{1'd0}, reg_}; // @[Memory.scala 23:14 Memory.scala 23:20 Memory.scala 22:18]
  assign io_out = {{1'd0}, reg_}; // @[Memory.scala 24:12]
  always @(posedge clock) begin
    reg_ <= _GEN_0[16:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_ = _RAND_0[16:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RandomHardware_1_16(
  input         clock,
  input  [18:0] io_in,
  output [17:0] io_out
);
  wire  RegE_000_clock; // @[RandomHardware_1_16.scala 14:26]
  wire [18:0] RegE_000_io_in; // @[RandomHardware_1_16.scala 14:26]
  wire [17:0] RegE_000_io_out; // @[RandomHardware_1_16.scala 14:26]
  RegE_3 RegE_000 ( // @[RandomHardware_1_16.scala 14:26]
    .clock(RegE_000_clock),
    .io_in(RegE_000_io_in),
    .io_out(RegE_000_io_out)
  );
  assign io_out = RegE_000_io_out; // @[RandomHardware_1_16.scala 17:10]
  assign RegE_000_clock = clock;
  assign RegE_000_io_in = io_in; // @[RandomHardware_1_16.scala 16:25]
endmodule
module ReduceOrMux(
  input  [15:0] io_in,
  output [5:0]  io_out
);
  wire [5:0] IN1 = io_in[15:10]; // @[Muxes.scala 110:27]
  wire [5:0] IN2 = io_in[9:4]; // @[Muxes.scala 111:27]
  wire [3:0] SEL = io_in[3:0]; // @[Muxes.scala 112:27]
  assign io_out = |SEL ? IN1 : IN2; // @[Muxes.scala 114:18]
endmodule
module RandomHardware_1_17(
  input  [15:0] io_in,
  output [5:0]  io_out
);
  wire [15:0] ReduceOrMux_000_io_in; // @[RandomHardware_1_17.scala 14:34]
  wire [5:0] ReduceOrMux_000_io_out; // @[RandomHardware_1_17.scala 14:34]
  ReduceOrMux ReduceOrMux_000 ( // @[RandomHardware_1_17.scala 14:34]
    .io_in(ReduceOrMux_000_io_in),
    .io_out(ReduceOrMux_000_io_out)
  );
  assign io_out = ReduceOrMux_000_io_out; // @[RandomHardware_1_17.scala 17:10]
  assign ReduceOrMux_000_io_in = io_in; // @[RandomHardware_1_17.scala 16:33]
endmodule
module ReduceXorMux_4(
  input  [39:0] io_in,
  output [14:0] io_out
);
  wire [14:0] IN1 = io_in[39:25]; // @[Muxes.scala 122:27]
  wire [14:0] IN2 = io_in[24:10]; // @[Muxes.scala 123:27]
  wire [9:0] SEL = io_in[9:0]; // @[Muxes.scala 124:27]
  assign io_out = ^SEL ? IN1 : IN2; // @[Muxes.scala 126:18]
endmodule
module RandomHardware_1_18(
  input         clock,
  input  [17:0] io_in,
  output [14:0] io_out
);
  wire  RandomHardware_000_clock; // @[RandomHardware_1_18.scala 15:42]
  wire [19:0] RandomHardware_000_io_in; // @[RandomHardware_1_18.scala 15:42]
  wire [7:0] RandomHardware_000_io_out; // @[RandomHardware_1_18.scala 15:42]
  wire [39:0] ReduceXorMux_001_io_in; // @[RandomHardware_1_18.scala 16:34]
  wire [14:0] ReduceXorMux_001_io_out; // @[RandomHardware_1_18.scala 16:34]
  RandomHardware_2_0 RandomHardware_000 ( // @[RandomHardware_1_18.scala 15:42]
    .clock(RandomHardware_000_clock),
    .io_in(RandomHardware_000_io_in),
    .io_out(RandomHardware_000_io_out)
  );
  ReduceXorMux_4 ReduceXorMux_001 ( // @[RandomHardware_1_18.scala 16:34]
    .io_in(ReduceXorMux_001_io_in),
    .io_out(ReduceXorMux_001_io_out)
  );
  assign io_out = ReduceXorMux_001_io_out; // @[RandomHardware_1_18.scala 19:10]
  assign RandomHardware_000_clock = clock;
  assign RandomHardware_000_io_in = {{2'd0}, io_in}; // @[RandomHardware_1_18.scala 18:33]
  assign ReduceXorMux_001_io_in = {{32'd0}, RandomHardware_000_io_out}; // @[RandomHardware_1_18.scala 13:24 RandomHardware_1_18.scala 21:18]
endmodule
module RandomHardware_1_19(
  input         clock,
  input  [19:0] io_in,
  output [7:0]  io_out
);
  wire  RandomHardware_000_clock; // @[RandomHardware_1_19.scala 14:42]
  wire [19:0] RandomHardware_000_io_in; // @[RandomHardware_1_19.scala 14:42]
  wire [7:0] RandomHardware_000_io_out; // @[RandomHardware_1_19.scala 14:42]
  RandomHardware_2_0 RandomHardware_000 ( // @[RandomHardware_1_19.scala 14:42]
    .clock(RandomHardware_000_clock),
    .io_in(RandomHardware_000_io_in),
    .io_out(RandomHardware_000_io_out)
  );
  assign io_out = RandomHardware_000_io_out; // @[RandomHardware_1_19.scala 17:10]
  assign RandomHardware_000_clock = clock;
  assign RandomHardware_000_io_in = io_in; // @[RandomHardware_1_19.scala 16:33]
endmodule
module RandomHardware_1_20(
  input  [19:0] io_in,
  output [7:0]  io_out
);
  wire [19:0] ReduceXorMux_000_io_in; // @[RandomHardware_1_20.scala 14:34]
  wire [7:0] ReduceXorMux_000_io_out; // @[RandomHardware_1_20.scala 14:34]
  ReduceXorMux ReduceXorMux_000 ( // @[RandomHardware_1_20.scala 14:34]
    .io_in(ReduceXorMux_000_io_in),
    .io_out(ReduceXorMux_000_io_out)
  );
  assign io_out = ReduceXorMux_000_io_out; // @[RandomHardware_1_20.scala 17:10]
  assign ReduceXorMux_000_io_in = io_in; // @[RandomHardware_1_20.scala 16:33]
endmodule
module SignExtendDouble_2(
  input  [5:0]  io_in,
  output [11:0] io_out
);
  wire [5:0] io_out_hi = io_in[5] ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  assign io_out = {io_out_hi,io_in}; // @[Cat.scala 30:58]
endmodule
module SignExtendDouble_3(
  input  [3:0] io_in,
  output [7:0] io_out
);
  wire [3:0] io_out_hi = io_in[3] ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  assign io_out = {io_out_hi,io_in}; // @[Cat.scala 30:58]
endmodule
module RandomHardware(
  input         clock,
  input         reset,
  input  [99:0] io_in,
  output [79:0] io_out
);
  wire [4:0] ShiftRight_000_io_in; // @[RandomHardware.scala 41:34]
  wire [4:0] ShiftRight_000_io_out; // @[RandomHardware.scala 41:34]
  wire [12:0] RandomHardware_001_io_in; // @[RandomHardware.scala 42:42]
  wire [12:0] RandomHardware_001_io_out; // @[RandomHardware.scala 42:42]
  wire  Accum_002_clock; // @[RandomHardware.scala 43:34]
  wire [7:0] Accum_002_io_in; // @[RandomHardware.scala 43:34]
  wire [7:0] Accum_002_io_out; // @[RandomHardware.scala 43:34]
  wire  RandomHardware_003_clock; // @[RandomHardware.scala 44:42]
  wire [15:0] RandomHardware_003_io_in; // @[RandomHardware.scala 44:42]
  wire [17:0] RandomHardware_003_io_out; // @[RandomHardware.scala 44:42]
  wire  RandomHardware_004_clock; // @[RandomHardware.scala 45:42]
  wire [36:0] RandomHardware_004_io_in; // @[RandomHardware.scala 45:42]
  wire [29:0] RandomHardware_004_io_out; // @[RandomHardware.scala 45:42]
  wire  ShiftRegister_005_clock; // @[RandomHardware.scala 46:42]
  wire [4:0] ShiftRegister_005_io_in; // @[RandomHardware.scala 46:42]
  wire [4:0] ShiftRegister_005_io_out; // @[RandomHardware.scala 46:42]
  wire  Reg_006_clock; // @[RandomHardware.scala 47:26]
  wire [7:0] Reg_006_io_in; // @[RandomHardware.scala 47:26]
  wire [7:0] Reg_006_io_out; // @[RandomHardware.scala 47:26]
  wire  RandomHardware_007_clock; // @[RandomHardware.scala 48:42]
  wire [20:0] RandomHardware_007_io_in; // @[RandomHardware.scala 48:42]
  wire [22:0] RandomHardware_007_io_out; // @[RandomHardware.scala 48:42]
  wire [15:0] RandomHardware_008_io_in; // @[RandomHardware.scala 49:42]
  wire [4:0] RandomHardware_008_io_out; // @[RandomHardware.scala 49:42]
  wire  ShiftRegister_009_clock; // @[RandomHardware.scala 50:42]
  wire [3:0] ShiftRegister_009_io_in; // @[RandomHardware.scala 50:42]
  wire [3:0] ShiftRegister_009_io_out; // @[RandomHardware.scala 50:42]
  wire  Accum_010_clock; // @[RandomHardware.scala 51:34]
  wire [5:0] Accum_010_io_in; // @[RandomHardware.scala 51:34]
  wire [5:0] Accum_010_io_out; // @[RandomHardware.scala 51:34]
  wire  RandomHardware_011_clock; // @[RandomHardware.scala 52:42]
  wire [15:0] RandomHardware_011_io_in; // @[RandomHardware.scala 52:42]
  wire [3:0] RandomHardware_011_io_out; // @[RandomHardware.scala 52:42]
  wire  RandomHardware_012_clock; // @[RandomHardware.scala 53:42]
  wire [11:0] RandomHardware_012_io_in; // @[RandomHardware.scala 53:42]
  wire [11:0] RandomHardware_012_io_out; // @[RandomHardware.scala 53:42]
  wire [18:0] RandomHardware_013_io_in; // @[RandomHardware.scala 54:42]
  wire [8:0] RandomHardware_013_io_out; // @[RandomHardware.scala 54:42]
  wire [5:0] Mul_014_io_in; // @[RandomHardware.scala 55:26]
  wire [5:0] Mul_014_io_out; // @[RandomHardware.scala 55:26]
  wire  Reg_015_clock; // @[RandomHardware.scala 56:26]
  wire [3:0] Reg_015_io_in; // @[RandomHardware.scala 56:26]
  wire [3:0] Reg_015_io_out; // @[RandomHardware.scala 56:26]
  wire  RandomHardware_016_clock; // @[RandomHardware.scala 57:42]
  wire [18:0] RandomHardware_016_io_in; // @[RandomHardware.scala 57:42]
  wire [17:0] RandomHardware_016_io_out; // @[RandomHardware.scala 57:42]
  wire [15:0] RandomHardware_017_io_in; // @[RandomHardware.scala 58:42]
  wire [5:0] RandomHardware_017_io_out; // @[RandomHardware.scala 58:42]
  wire  RandomHardware_018_clock; // @[RandomHardware.scala 59:42]
  wire [17:0] RandomHardware_018_io_in; // @[RandomHardware.scala 59:42]
  wire [14:0] RandomHardware_018_io_out; // @[RandomHardware.scala 59:42]
  wire  RandomHardware_019_clock; // @[RandomHardware.scala 60:42]
  wire [19:0] RandomHardware_019_io_in; // @[RandomHardware.scala 60:42]
  wire [7:0] RandomHardware_019_io_out; // @[RandomHardware.scala 60:42]
  wire [19:0] RandomHardware_020_io_in; // @[RandomHardware.scala 61:42]
  wire [7:0] RandomHardware_020_io_out; // @[RandomHardware.scala 61:42]
  wire  ShiftRegister_021_clock; // @[RandomHardware.scala 62:42]
  wire [4:0] ShiftRegister_021_io_in; // @[RandomHardware.scala 62:42]
  wire [4:0] ShiftRegister_021_io_out; // @[RandomHardware.scala 62:42]
  wire [5:0] SignExtendDouble_022_io_in; // @[RandomHardware.scala 63:42]
  wire [11:0] SignExtendDouble_022_io_out; // @[RandomHardware.scala 63:42]
  wire [3:0] SignExtendDouble_023_io_in; // @[RandomHardware.scala 64:42]
  wire [7:0] SignExtendDouble_023_io_out; // @[RandomHardware.scala 64:42]
  wire  Accum_024_clock; // @[RandomHardware.scala 65:34]
  wire [5:0] Accum_024_io_in; // @[RandomHardware.scala 65:34]
  wire [5:0] Accum_024_io_out; // @[RandomHardware.scala 65:34]
  wire [31:0] io_out_lo = {Reg_006_io_out,Mul_014_io_out,RandomHardware_016_io_out}; // @[Cat.scala 30:58]
  wire [47:0] io_out_hi = {ShiftRight_000_io_out,RandomHardware_001_io_out,RandomHardware_004_io_out}; // @[Cat.scala 30:58]
  wire [3:0] wire_004 = RandomHardware_011_io_out; // @[RandomHardware.scala 17:24 RandomHardware.scala 108:18]
  wire [11:0] wire_005 = RandomHardware_012_io_out; // @[RandomHardware.scala 18:24 RandomHardware.scala 111:18]
  wire [8:0] wire_011 = RandomHardware_013_io_out; // @[RandomHardware.scala 24:24 RandomHardware.scala 93:18]
  wire [11:0] wire_012 = SignExtendDouble_022_io_out; // @[RandomHardware.scala 25:24 RandomHardware.scala 102:18]
  wire [7:0] wire_015 = Accum_002_io_out; // @[RandomHardware.scala 28:24 RandomHardware.scala 77:18]
  wire [4:0] wire_016 = ShiftRegister_021_io_out; // @[RandomHardware.scala 29:24 RandomHardware.scala 100:18]
  wire [12:0] RandomHardware_013_io_in_hi = {wire_015,wire_016}; // @[Cat.scala 30:58]
  wire [5:0] wire_017 = Accum_024_io_out; // @[RandomHardware.scala 30:24 RandomHardware.scala 106:18]
  wire [7:0] wire_002 = SignExtendDouble_023_io_out; // @[RandomHardware.scala 15:24 RandomHardware.scala 104:18]
  wire [22:0] wire_006 = RandomHardware_007_io_out; // @[RandomHardware.scala 19:24 RandomHardware.scala 84:18]
  wire [5:0] wire_007 = Accum_010_io_out; // @[RandomHardware.scala 20:24 RandomHardware.scala 88:18]
  wire [28:0] RandomHardware_004_io_in_hi = {wire_006,wire_007}; // @[Cat.scala 30:58]
  wire [7:0] wire_008 = RandomHardware_019_io_out; // @[RandomHardware.scala 21:24 RandomHardware.scala 113:18]
  wire [14:0] wire_021 = RandomHardware_018_io_out; // @[RandomHardware.scala 34:24 RandomHardware.scala 97:18]
  ShiftRight ShiftRight_000 ( // @[RandomHardware.scala 41:34]
    .io_in(ShiftRight_000_io_in),
    .io_out(ShiftRight_000_io_out)
  );
  RandomHardware_1_1 RandomHardware_001 ( // @[RandomHardware.scala 42:42]
    .io_in(RandomHardware_001_io_in),
    .io_out(RandomHardware_001_io_out)
  );
  Accum Accum_002 ( // @[RandomHardware.scala 43:34]
    .clock(Accum_002_clock),
    .io_in(Accum_002_io_in),
    .io_out(Accum_002_io_out)
  );
  RandomHardware_1_3 RandomHardware_003 ( // @[RandomHardware.scala 44:42]
    .clock(RandomHardware_003_clock),
    .io_in(RandomHardware_003_io_in),
    .io_out(RandomHardware_003_io_out)
  );
  RandomHardware_1_4 RandomHardware_004 ( // @[RandomHardware.scala 45:42]
    .clock(RandomHardware_004_clock),
    .io_in(RandomHardware_004_io_in),
    .io_out(RandomHardware_004_io_out)
  );
  ShiftRegister ShiftRegister_005 ( // @[RandomHardware.scala 46:42]
    .clock(ShiftRegister_005_clock),
    .io_in(ShiftRegister_005_io_in),
    .io_out(ShiftRegister_005_io_out)
  );
  Reg_1 Reg_006 ( // @[RandomHardware.scala 47:26]
    .clock(Reg_006_clock),
    .io_in(Reg_006_io_in),
    .io_out(Reg_006_io_out)
  );
  RandomHardware_1_7 RandomHardware_007 ( // @[RandomHardware.scala 48:42]
    .clock(RandomHardware_007_clock),
    .io_in(RandomHardware_007_io_in),
    .io_out(RandomHardware_007_io_out)
  );
  RandomHardware_1_8 RandomHardware_008 ( // @[RandomHardware.scala 49:42]
    .io_in(RandomHardware_008_io_in),
    .io_out(RandomHardware_008_io_out)
  );
  ShiftRegister_1 ShiftRegister_009 ( // @[RandomHardware.scala 50:42]
    .clock(ShiftRegister_009_clock),
    .io_in(ShiftRegister_009_io_in),
    .io_out(ShiftRegister_009_io_out)
  );
  Accum_2 Accum_010 ( // @[RandomHardware.scala 51:34]
    .clock(Accum_010_clock),
    .io_in(Accum_010_io_in),
    .io_out(Accum_010_io_out)
  );
  RandomHardware_1_11 RandomHardware_011 ( // @[RandomHardware.scala 52:42]
    .clock(RandomHardware_011_clock),
    .io_in(RandomHardware_011_io_in),
    .io_out(RandomHardware_011_io_out)
  );
  RandomHardware_1_12 RandomHardware_012 ( // @[RandomHardware.scala 53:42]
    .clock(RandomHardware_012_clock),
    .io_in(RandomHardware_012_io_in),
    .io_out(RandomHardware_012_io_out)
  );
  RandomHardware_1_13 RandomHardware_013 ( // @[RandomHardware.scala 54:42]
    .io_in(RandomHardware_013_io_in),
    .io_out(RandomHardware_013_io_out)
  );
  Mul Mul_014 ( // @[RandomHardware.scala 55:26]
    .io_in(Mul_014_io_in),
    .io_out(Mul_014_io_out)
  );
  Reg_2 Reg_015 ( // @[RandomHardware.scala 56:26]
    .clock(Reg_015_clock),
    .io_in(Reg_015_io_in),
    .io_out(Reg_015_io_out)
  );
  RandomHardware_1_16 RandomHardware_016 ( // @[RandomHardware.scala 57:42]
    .clock(RandomHardware_016_clock),
    .io_in(RandomHardware_016_io_in),
    .io_out(RandomHardware_016_io_out)
  );
  RandomHardware_1_17 RandomHardware_017 ( // @[RandomHardware.scala 58:42]
    .io_in(RandomHardware_017_io_in),
    .io_out(RandomHardware_017_io_out)
  );
  RandomHardware_1_18 RandomHardware_018 ( // @[RandomHardware.scala 59:42]
    .clock(RandomHardware_018_clock),
    .io_in(RandomHardware_018_io_in),
    .io_out(RandomHardware_018_io_out)
  );
  RandomHardware_1_19 RandomHardware_019 ( // @[RandomHardware.scala 60:42]
    .clock(RandomHardware_019_clock),
    .io_in(RandomHardware_019_io_in),
    .io_out(RandomHardware_019_io_out)
  );
  RandomHardware_1_20 RandomHardware_020 ( // @[RandomHardware.scala 61:42]
    .io_in(RandomHardware_020_io_in),
    .io_out(RandomHardware_020_io_out)
  );
  ShiftRegister ShiftRegister_021 ( // @[RandomHardware.scala 62:42]
    .clock(ShiftRegister_021_clock),
    .io_in(ShiftRegister_021_io_in),
    .io_out(ShiftRegister_021_io_out)
  );
  SignExtendDouble_2 SignExtendDouble_022 ( // @[RandomHardware.scala 63:42]
    .io_in(SignExtendDouble_022_io_in),
    .io_out(SignExtendDouble_022_io_out)
  );
  SignExtendDouble_3 SignExtendDouble_023 ( // @[RandomHardware.scala 64:42]
    .io_in(SignExtendDouble_023_io_in),
    .io_out(SignExtendDouble_023_io_out)
  );
  Accum_2 Accum_024 ( // @[RandomHardware.scala 65:34]
    .clock(Accum_024_clock),
    .io_in(Accum_024_io_in),
    .io_out(Accum_024_io_out)
  );
  assign io_out = {io_out_hi,io_out_lo}; // @[Cat.scala 30:58]
  assign ShiftRight_000_io_in = ShiftRegister_005_io_out; // @[RandomHardware.scala 13:24 RandomHardware.scala 81:18]
  assign RandomHardware_001_io_in = {wire_016,wire_002}; // @[Cat.scala 30:58]
  assign Accum_002_clock = clock;
  assign Accum_002_io_in = RandomHardware_020_io_out; // @[RandomHardware.scala 16:24 RandomHardware.scala 114:18]
  assign RandomHardware_003_clock = clock;
  assign RandomHardware_003_io_in = {wire_004,wire_005}; // @[Cat.scala 30:58]
  assign RandomHardware_004_clock = clock;
  assign RandomHardware_004_io_in = {RandomHardware_004_io_in_hi,wire_008}; // @[Cat.scala 30:58]
  assign ShiftRegister_005_clock = clock;
  assign ShiftRegister_005_io_in = RandomHardware_008_io_out; // @[RandomHardware.scala 22:24 RandomHardware.scala 107:18]
  assign Reg_006_clock = clock;
  assign Reg_006_io_in = Accum_002_io_out; // @[RandomHardware.scala 23:24 RandomHardware.scala 76:18]
  assign RandomHardware_007_clock = clock;
  assign RandomHardware_007_io_in = {wire_011,wire_012}; // @[Cat.scala 30:58]
  assign RandomHardware_008_io_in = io_in[15:0]; // @[RandomHardware.scala 67:41]
  assign ShiftRegister_009_clock = clock;
  assign ShiftRegister_009_io_in = Reg_015_io_out; // @[RandomHardware.scala 26:24 RandomHardware.scala 95:18]
  assign Accum_010_clock = clock;
  assign Accum_010_io_in = RandomHardware_017_io_out; // @[RandomHardware.scala 27:24 RandomHardware.scala 112:18]
  assign RandomHardware_011_clock = clock;
  assign RandomHardware_011_io_in = io_in[99:84]; // @[RandomHardware.scala 68:41]
  assign RandomHardware_012_clock = clock;
  assign RandomHardware_012_io_in = io_in[99:88]; // @[RandomHardware.scala 69:41]
  assign RandomHardware_013_io_in = {RandomHardware_013_io_in_hi,wire_017}; // @[Cat.scala 30:58]
  assign Mul_014_io_in = Accum_010_io_out; // @[RandomHardware.scala 31:24 RandomHardware.scala 89:18]
  assign Reg_015_clock = clock;
  assign Reg_015_io_in = RandomHardware_011_io_out; // @[RandomHardware.scala 32:24 RandomHardware.scala 109:18]
  assign RandomHardware_016_clock = clock;
  assign RandomHardware_016_io_in = {wire_004,wire_021}; // @[Cat.scala 30:58]
  assign RandomHardware_017_io_in = io_in[15:0]; // @[RandomHardware.scala 70:41]
  assign RandomHardware_018_clock = clock;
  assign RandomHardware_018_io_in = RandomHardware_003_io_out; // @[RandomHardware.scala 35:24 RandomHardware.scala 79:18]
  assign RandomHardware_019_clock = clock;
  assign RandomHardware_019_io_in = io_in[99:80]; // @[RandomHardware.scala 71:41]
  assign RandomHardware_020_io_in = io_in[19:0]; // @[RandomHardware.scala 72:41]
  assign ShiftRegister_021_clock = clock;
  assign ShiftRegister_021_io_in = ShiftRegister_005_io_out; // @[RandomHardware.scala 36:24 RandomHardware.scala 82:18]
  assign SignExtendDouble_022_io_in = Accum_010_io_out; // @[RandomHardware.scala 37:24 RandomHardware.scala 90:18]
  assign SignExtendDouble_023_io_in = ShiftRegister_009_io_out; // @[RandomHardware.scala 38:24 RandomHardware.scala 86:18]
  assign Accum_024_clock = clock;
  assign Accum_024_io_in = Accum_010_io_out; // @[RandomHardware.scala 39:24 RandomHardware.scala 91:18]
endmodule
