module ComputeAdd(
  input  [25:0] io_in1,
  input  [25:0] io_in2,
  output [52:0] io_out
);
  wire [25:0] _io_out_T_1 = io_in1 + io_in2; // @[Arithmetics.scala 13:22]
  assign io_out = {{27'd0}, _io_out_T_1}; // @[Arithmetics.scala 13:22]
endmodule
module ComputeAdd_1(
  input        io_in1,
  input        io_in2,
  output [1:0] io_out
);
  wire  _io_out_T_1 = io_in1 + io_in2; // @[Arithmetics.scala 13:22]
  assign io_out = {{1'd0}, _io_out_T_1}; // @[Arithmetics.scala 13:22]
endmodule
module ComputeAdd_2(
  input  [1:0] io_in1,
  input  [1:0] io_in2,
  output [4:0] io_out
);
  wire [1:0] _io_out_T_1 = io_in1 + io_in2; // @[Arithmetics.scala 13:22]
  assign io_out = {{3'd0}, _io_out_T_1}; // @[Arithmetics.scala 13:22]
endmodule
module ComputeAdd_3(
  input  [2:0] io_in1,
  input  [2:0] io_in2,
  output [6:0] io_out
);
  wire [2:0] _io_out_T_1 = io_in1 + io_in2; // @[Arithmetics.scala 13:22]
  assign io_out = {{4'd0}, _io_out_T_1}; // @[Arithmetics.scala 13:22]
endmodule
module ComputeAdd_5(
  input  [7:0]  io_in1,
  input  [7:0]  io_in2,
  output [15:0] io_out
);
  wire [7:0] _io_out_T_1 = io_in1 + io_in2; // @[Arithmetics.scala 13:22]
  assign io_out = {{8'd0}, _io_out_T_1}; // @[Arithmetics.scala 13:22]
endmodule
module ComputeAdd_7(
  input  [8:0]  io_in1,
  input  [8:0]  io_in2,
  output [17:0] io_out
);
  wire [8:0] _io_out_T_1 = io_in1 + io_in2; // @[Arithmetics.scala 13:22]
  assign io_out = {{9'd0}, _io_out_T_1}; // @[Arithmetics.scala 13:22]
endmodule
module ComputeAdd_8(
  input  [6:0]  io_in1,
  input  [6:0]  io_in2,
  output [13:0] io_out
);
  wire [6:0] _io_out_T_1 = io_in1 + io_in2; // @[Arithmetics.scala 13:22]
  assign io_out = {{7'd0}, _io_out_T_1}; // @[Arithmetics.scala 13:22]
endmodule
module ComputeAdd_9(
  input  [3:0] io_in1,
  input  [3:0] io_in2,
  output [7:0] io_out
);
  wire [3:0] _io_out_T_1 = io_in1 + io_in2; // @[Arithmetics.scala 13:22]
  assign io_out = {{4'd0}, _io_out_T_1}; // @[Arithmetics.scala 13:22]
endmodule
module ComputeAdd_10(
  input  [4:0] io_in1,
  input  [4:0] io_in2,
  output [9:0] io_out
);
  wire [4:0] _io_out_T_1 = io_in1 + io_in2; // @[Arithmetics.scala 13:22]
  assign io_out = {{5'd0}, _io_out_T_1}; // @[Arithmetics.scala 13:22]
endmodule
module ComputeAdd_17(
  input  [5:0]  io_in1,
  input  [5:0]  io_in2,
  output [11:0] io_out
);
  wire [5:0] _io_out_T_1 = io_in1 + io_in2; // @[Arithmetics.scala 13:22]
  assign io_out = {{6'd0}, _io_out_T_1}; // @[Arithmetics.scala 13:22]
endmodule
module ComputeAdd_18(
  input  [1:0] io_in1,
  input  [1:0] io_in2,
  output [3:0] io_out
);
  wire [1:0] _io_out_T_1 = io_in1 + io_in2; // @[Arithmetics.scala 13:22]
  assign io_out = {{2'd0}, _io_out_T_1}; // @[Arithmetics.scala 13:22]
endmodule
module RandomHardware(
  input         clock,
  input         reset,
  input  [97:0] io_in,
  output [95:0] io_out
);
  wire [25:0] Comp_Adder_000_io_in1; // @[RandomHardware.scala 34:34]
  wire [25:0] Comp_Adder_000_io_in2; // @[RandomHardware.scala 34:34]
  wire [52:0] Comp_Adder_000_io_out; // @[RandomHardware.scala 34:34]
  wire  Comp_Adder_001_io_in1; // @[RandomHardware.scala 35:34]
  wire  Comp_Adder_001_io_in2; // @[RandomHardware.scala 35:34]
  wire [1:0] Comp_Adder_001_io_out; // @[RandomHardware.scala 35:34]
  wire [1:0] Comp_Adder_002_io_in1; // @[RandomHardware.scala 36:34]
  wire [1:0] Comp_Adder_002_io_in2; // @[RandomHardware.scala 36:34]
  wire [4:0] Comp_Adder_002_io_out; // @[RandomHardware.scala 36:34]
  wire [2:0] Comp_Adder_003_io_in1; // @[RandomHardware.scala 37:34]
  wire [2:0] Comp_Adder_003_io_in2; // @[RandomHardware.scala 37:34]
  wire [6:0] Comp_Adder_003_io_out; // @[RandomHardware.scala 37:34]
  wire  Comp_Adder_004_io_in1; // @[RandomHardware.scala 38:34]
  wire  Comp_Adder_004_io_in2; // @[RandomHardware.scala 38:34]
  wire [1:0] Comp_Adder_004_io_out; // @[RandomHardware.scala 38:34]
  wire [7:0] Comp_Adder_005_io_in1; // @[RandomHardware.scala 39:34]
  wire [7:0] Comp_Adder_005_io_in2; // @[RandomHardware.scala 39:34]
  wire [15:0] Comp_Adder_005_io_out; // @[RandomHardware.scala 39:34]
  wire  Comp_Adder_006_io_in1; // @[RandomHardware.scala 40:34]
  wire  Comp_Adder_006_io_in2; // @[RandomHardware.scala 40:34]
  wire [1:0] Comp_Adder_006_io_out; // @[RandomHardware.scala 40:34]
  wire [8:0] Comp_Adder_007_io_in1; // @[RandomHardware.scala 41:34]
  wire [8:0] Comp_Adder_007_io_in2; // @[RandomHardware.scala 41:34]
  wire [17:0] Comp_Adder_007_io_out; // @[RandomHardware.scala 41:34]
  wire [6:0] Comp_Adder_008_io_in1; // @[RandomHardware.scala 42:34]
  wire [6:0] Comp_Adder_008_io_in2; // @[RandomHardware.scala 42:34]
  wire [13:0] Comp_Adder_008_io_out; // @[RandomHardware.scala 42:34]
  wire [3:0] Comp_Adder_009_io_in1; // @[RandomHardware.scala 43:34]
  wire [3:0] Comp_Adder_009_io_in2; // @[RandomHardware.scala 43:34]
  wire [7:0] Comp_Adder_009_io_out; // @[RandomHardware.scala 43:34]
  wire [4:0] Comp_Adder_010_io_in1; // @[RandomHardware.scala 44:34]
  wire [4:0] Comp_Adder_010_io_in2; // @[RandomHardware.scala 44:34]
  wire [9:0] Comp_Adder_010_io_out; // @[RandomHardware.scala 44:34]
  wire [3:0] Comp_Adder_011_io_in1; // @[RandomHardware.scala 45:34]
  wire [3:0] Comp_Adder_011_io_in2; // @[RandomHardware.scala 45:34]
  wire [7:0] Comp_Adder_011_io_out; // @[RandomHardware.scala 45:34]
  wire [6:0] Comp_Adder_012_io_in1; // @[RandomHardware.scala 46:34]
  wire [6:0] Comp_Adder_012_io_in2; // @[RandomHardware.scala 46:34]
  wire [13:0] Comp_Adder_012_io_out; // @[RandomHardware.scala 46:34]
  wire [1:0] Comp_Adder_013_io_in1; // @[RandomHardware.scala 47:34]
  wire [1:0] Comp_Adder_013_io_in2; // @[RandomHardware.scala 47:34]
  wire [4:0] Comp_Adder_013_io_out; // @[RandomHardware.scala 47:34]
  wire [2:0] Comp_Adder_014_io_in1; // @[RandomHardware.scala 48:34]
  wire [2:0] Comp_Adder_014_io_in2; // @[RandomHardware.scala 48:34]
  wire [6:0] Comp_Adder_014_io_out; // @[RandomHardware.scala 48:34]
  wire [4:0] Comp_Adder_015_io_in1; // @[RandomHardware.scala 49:34]
  wire [4:0] Comp_Adder_015_io_in2; // @[RandomHardware.scala 49:34]
  wire [9:0] Comp_Adder_015_io_out; // @[RandomHardware.scala 49:34]
  wire [2:0] Comp_Adder_016_io_in1; // @[RandomHardware.scala 50:34]
  wire [2:0] Comp_Adder_016_io_in2; // @[RandomHardware.scala 50:34]
  wire [6:0] Comp_Adder_016_io_out; // @[RandomHardware.scala 50:34]
  wire [5:0] Comp_Adder_017_io_in1; // @[RandomHardware.scala 51:34]
  wire [5:0] Comp_Adder_017_io_in2; // @[RandomHardware.scala 51:34]
  wire [11:0] Comp_Adder_017_io_out; // @[RandomHardware.scala 51:34]
  wire [1:0] Comp_Adder_018_io_in1; // @[RandomHardware.scala 52:34]
  wire [1:0] Comp_Adder_018_io_in2; // @[RandomHardware.scala 52:34]
  wire [3:0] Comp_Adder_018_io_out; // @[RandomHardware.scala 52:34]
  wire [6:0] Comp_Adder_019_io_in1; // @[RandomHardware.scala 53:34]
  wire [6:0] Comp_Adder_019_io_in2; // @[RandomHardware.scala 53:34]
  wire [13:0] Comp_Adder_019_io_out; // @[RandomHardware.scala 53:34]
  wire [3:0] Comp_Adder_020_io_in1; // @[RandomHardware.scala 54:34]
  wire [3:0] Comp_Adder_020_io_in2; // @[RandomHardware.scala 54:34]
  wire [7:0] Comp_Adder_020_io_out; // @[RandomHardware.scala 54:34]
  wire [17:0] io_out_lo = {Comp_Adder_014_io_out,Comp_Adder_016_io_out,Comp_Adder_018_io_out}; // @[Cat.scala 30:58]
  wire [77:0] io_out_hi = {Comp_Adder_000_io_out,Comp_Adder_004_io_out,Comp_Adder_007_io_out,Comp_Adder_013_io_out}; // @[Cat.scala 30:58]
  wire [1:0] temp_vertex_001 = Comp_Adder_003_io_out[1:0]; // @[RandomHardware.scala 85:43]
  wire [1:0] temp_vertex_006 = Comp_Adder_001_io_out; // @[RandomHardware.scala 77:43]
  wire [4:0] temp_vertex_002 = Comp_Adder_010_io_out[4:0]; // @[RandomHardware.scala 104:43]
  wire [4:0] wire_019 = Comp_Adder_002_io_out; // @[RandomHardware.scala 81:43]
  wire [6:0] temp_vertex_003 = Comp_Adder_019_io_out[6:0]; // @[RandomHardware.scala 111:43]
  wire [1:0] temp_vertex_004 = Comp_Adder_003_io_out[3:2]; // @[RandomHardware.scala 86:43]
  wire [2:0] wire_020 = Comp_Adder_003_io_out[6:4]; // @[RandomHardware.scala 87:43]
  wire [1:0] wire_010 = Comp_Adder_006_io_out; // @[RandomHardware.scala 91:43]
  wire [7:0] temp_vertex_009 = Comp_Adder_011_io_out; // @[RandomHardware.scala 106:43]
  wire [3:0] wire_012 = Comp_Adder_009_io_out[3:0]; // @[RandomHardware.scala 95:43]
  wire [3:0] temp_vertex_018 = Comp_Adder_009_io_out[7:4]; // @[RandomHardware.scala 96:43]
  wire [7:0] temp_vertex_020 = {wire_019,wire_020}; // @[Cat.scala 30:58]
  wire [7:0] wire_004 = Comp_Adder_020_io_out; // @[RandomHardware.scala 100:43]
  wire [15:0] wire_000 = Comp_Adder_005_io_out; // @[RandomHardware.scala 101:43]
  wire [6:0] wire_011 = Comp_Adder_008_io_out[6:0]; // @[RandomHardware.scala 102:43]
  wire [6:0] temp_vertex_014 = Comp_Adder_008_io_out[13:7]; // @[RandomHardware.scala 103:43]
  wire [4:0] temp_vertex_013 = Comp_Adder_010_io_out[9:5]; // @[RandomHardware.scala 105:43]
  wire [6:0] wire_001 = Comp_Adder_012_io_out[6:0]; // @[RandomHardware.scala 107:43]
  wire [6:0] temp_vertex_016 = Comp_Adder_012_io_out[13:7]; // @[RandomHardware.scala 108:43]
  wire [9:0] wire_002 = Comp_Adder_015_io_out; // @[RandomHardware.scala 109:43]
  wire [11:0] wire_003 = Comp_Adder_017_io_out; // @[RandomHardware.scala 110:43]
  wire [6:0] wire_013 = Comp_Adder_019_io_out[13:7]; // @[RandomHardware.scala 112:43]
  wire [52:0] temp_vertex_000 = {wire_000,wire_001,wire_002,wire_003,wire_004}; // @[Cat.scala 30:58]
  wire [19:0] temp_vertex_007 = {wire_010,wire_011,wire_012,wire_013}; // @[Cat.scala 30:58]
  ComputeAdd Comp_Adder_000 ( // @[RandomHardware.scala 34:34]
    .io_in1(Comp_Adder_000_io_in1),
    .io_in2(Comp_Adder_000_io_in2),
    .io_out(Comp_Adder_000_io_out)
  );
  ComputeAdd_1 Comp_Adder_001 ( // @[RandomHardware.scala 35:34]
    .io_in1(Comp_Adder_001_io_in1),
    .io_in2(Comp_Adder_001_io_in2),
    .io_out(Comp_Adder_001_io_out)
  );
  ComputeAdd_2 Comp_Adder_002 ( // @[RandomHardware.scala 36:34]
    .io_in1(Comp_Adder_002_io_in1),
    .io_in2(Comp_Adder_002_io_in2),
    .io_out(Comp_Adder_002_io_out)
  );
  ComputeAdd_3 Comp_Adder_003 ( // @[RandomHardware.scala 37:34]
    .io_in1(Comp_Adder_003_io_in1),
    .io_in2(Comp_Adder_003_io_in2),
    .io_out(Comp_Adder_003_io_out)
  );
  ComputeAdd_1 Comp_Adder_004 ( // @[RandomHardware.scala 38:34]
    .io_in1(Comp_Adder_004_io_in1),
    .io_in2(Comp_Adder_004_io_in2),
    .io_out(Comp_Adder_004_io_out)
  );
  ComputeAdd_5 Comp_Adder_005 ( // @[RandomHardware.scala 39:34]
    .io_in1(Comp_Adder_005_io_in1),
    .io_in2(Comp_Adder_005_io_in2),
    .io_out(Comp_Adder_005_io_out)
  );
  ComputeAdd_1 Comp_Adder_006 ( // @[RandomHardware.scala 40:34]
    .io_in1(Comp_Adder_006_io_in1),
    .io_in2(Comp_Adder_006_io_in2),
    .io_out(Comp_Adder_006_io_out)
  );
  ComputeAdd_7 Comp_Adder_007 ( // @[RandomHardware.scala 41:34]
    .io_in1(Comp_Adder_007_io_in1),
    .io_in2(Comp_Adder_007_io_in2),
    .io_out(Comp_Adder_007_io_out)
  );
  ComputeAdd_8 Comp_Adder_008 ( // @[RandomHardware.scala 42:34]
    .io_in1(Comp_Adder_008_io_in1),
    .io_in2(Comp_Adder_008_io_in2),
    .io_out(Comp_Adder_008_io_out)
  );
  ComputeAdd_9 Comp_Adder_009 ( // @[RandomHardware.scala 43:34]
    .io_in1(Comp_Adder_009_io_in1),
    .io_in2(Comp_Adder_009_io_in2),
    .io_out(Comp_Adder_009_io_out)
  );
  ComputeAdd_10 Comp_Adder_010 ( // @[RandomHardware.scala 44:34]
    .io_in1(Comp_Adder_010_io_in1),
    .io_in2(Comp_Adder_010_io_in2),
    .io_out(Comp_Adder_010_io_out)
  );
  ComputeAdd_9 Comp_Adder_011 ( // @[RandomHardware.scala 45:34]
    .io_in1(Comp_Adder_011_io_in1),
    .io_in2(Comp_Adder_011_io_in2),
    .io_out(Comp_Adder_011_io_out)
  );
  ComputeAdd_8 Comp_Adder_012 ( // @[RandomHardware.scala 46:34]
    .io_in1(Comp_Adder_012_io_in1),
    .io_in2(Comp_Adder_012_io_in2),
    .io_out(Comp_Adder_012_io_out)
  );
  ComputeAdd_2 Comp_Adder_013 ( // @[RandomHardware.scala 47:34]
    .io_in1(Comp_Adder_013_io_in1),
    .io_in2(Comp_Adder_013_io_in2),
    .io_out(Comp_Adder_013_io_out)
  );
  ComputeAdd_3 Comp_Adder_014 ( // @[RandomHardware.scala 48:34]
    .io_in1(Comp_Adder_014_io_in1),
    .io_in2(Comp_Adder_014_io_in2),
    .io_out(Comp_Adder_014_io_out)
  );
  ComputeAdd_10 Comp_Adder_015 ( // @[RandomHardware.scala 49:34]
    .io_in1(Comp_Adder_015_io_in1),
    .io_in2(Comp_Adder_015_io_in2),
    .io_out(Comp_Adder_015_io_out)
  );
  ComputeAdd_3 Comp_Adder_016 ( // @[RandomHardware.scala 50:34]
    .io_in1(Comp_Adder_016_io_in1),
    .io_in2(Comp_Adder_016_io_in2),
    .io_out(Comp_Adder_016_io_out)
  );
  ComputeAdd_17 Comp_Adder_017 ( // @[RandomHardware.scala 51:34]
    .io_in1(Comp_Adder_017_io_in1),
    .io_in2(Comp_Adder_017_io_in2),
    .io_out(Comp_Adder_017_io_out)
  );
  ComputeAdd_18 Comp_Adder_018 ( // @[RandomHardware.scala 52:34]
    .io_in1(Comp_Adder_018_io_in1),
    .io_in2(Comp_Adder_018_io_in2),
    .io_out(Comp_Adder_018_io_out)
  );
  ComputeAdd_8 Comp_Adder_019 ( // @[RandomHardware.scala 53:34]
    .io_in1(Comp_Adder_019_io_in1),
    .io_in2(Comp_Adder_019_io_in2),
    .io_out(Comp_Adder_019_io_out)
  );
  ComputeAdd_9 Comp_Adder_020 ( // @[RandomHardware.scala 54:34]
    .io_in1(Comp_Adder_020_io_in1),
    .io_in2(Comp_Adder_020_io_in2),
    .io_out(Comp_Adder_020_io_out)
  );
  assign io_out = {io_out_hi,io_out_lo}; // @[Cat.scala 30:58]
  assign Comp_Adder_000_io_in1 = temp_vertex_000[25:0]; // @[RandomHardware.scala 114:51]
  assign Comp_Adder_000_io_in2 = temp_vertex_000[51:26]; // @[RandomHardware.scala 115:33]
  assign Comp_Adder_001_io_in1 = temp_vertex_001[0]; // @[RandomHardware.scala 75:51]
  assign Comp_Adder_001_io_in2 = temp_vertex_001[1]; // @[RandomHardware.scala 76:51]
  assign Comp_Adder_002_io_in1 = temp_vertex_002[1:0]; // @[RandomHardware.scala 79:51]
  assign Comp_Adder_002_io_in2 = temp_vertex_002[3:2]; // @[RandomHardware.scala 80:33]
  assign Comp_Adder_003_io_in1 = temp_vertex_003[2:0]; // @[RandomHardware.scala 83:51]
  assign Comp_Adder_003_io_in2 = temp_vertex_003[5:3]; // @[RandomHardware.scala 84:33]
  assign Comp_Adder_004_io_in1 = temp_vertex_004[0]; // @[RandomHardware.scala 117:51]
  assign Comp_Adder_004_io_in2 = temp_vertex_004[1]; // @[RandomHardware.scala 118:51]
  assign Comp_Adder_005_io_in1 = io_in[7:0]; // @[RandomHardware.scala 56:41]
  assign Comp_Adder_005_io_in2 = io_in[15:8]; // @[RandomHardware.scala 57:41]
  assign Comp_Adder_006_io_in1 = temp_vertex_006[0]; // @[RandomHardware.scala 89:51]
  assign Comp_Adder_006_io_in2 = temp_vertex_006[1]; // @[RandomHardware.scala 90:51]
  assign Comp_Adder_007_io_in1 = temp_vertex_007[8:0]; // @[RandomHardware.scala 120:51]
  assign Comp_Adder_007_io_in2 = temp_vertex_007[17:9]; // @[RandomHardware.scala 121:51]
  assign Comp_Adder_008_io_in1 = io_in[22:16]; // @[RandomHardware.scala 58:41]
  assign Comp_Adder_008_io_in2 = io_in[29:23]; // @[RandomHardware.scala 59:41]
  assign Comp_Adder_009_io_in1 = temp_vertex_009[3:0]; // @[RandomHardware.scala 93:51]
  assign Comp_Adder_009_io_in2 = temp_vertex_009[7:4]; // @[RandomHardware.scala 94:51]
  assign Comp_Adder_010_io_in1 = io_in[34:30]; // @[RandomHardware.scala 60:41]
  assign Comp_Adder_010_io_in2 = io_in[39:35]; // @[RandomHardware.scala 61:41]
  assign Comp_Adder_011_io_in1 = io_in[43:40]; // @[RandomHardware.scala 62:41]
  assign Comp_Adder_011_io_in2 = io_in[47:44]; // @[RandomHardware.scala 63:41]
  assign Comp_Adder_012_io_in1 = io_in[54:48]; // @[RandomHardware.scala 64:41]
  assign Comp_Adder_012_io_in2 = io_in[61:55]; // @[RandomHardware.scala 65:41]
  assign Comp_Adder_013_io_in1 = temp_vertex_013[1:0]; // @[RandomHardware.scala 123:51]
  assign Comp_Adder_013_io_in2 = temp_vertex_013[3:2]; // @[RandomHardware.scala 124:33]
  assign Comp_Adder_014_io_in1 = temp_vertex_014[2:0]; // @[RandomHardware.scala 126:51]
  assign Comp_Adder_014_io_in2 = temp_vertex_014[5:3]; // @[RandomHardware.scala 127:33]
  assign Comp_Adder_015_io_in1 = io_in[66:62]; // @[RandomHardware.scala 66:41]
  assign Comp_Adder_015_io_in2 = io_in[71:67]; // @[RandomHardware.scala 67:41]
  assign Comp_Adder_016_io_in1 = temp_vertex_016[2:0]; // @[RandomHardware.scala 129:51]
  assign Comp_Adder_016_io_in2 = temp_vertex_016[5:3]; // @[RandomHardware.scala 130:33]
  assign Comp_Adder_017_io_in1 = io_in[77:72]; // @[RandomHardware.scala 68:41]
  assign Comp_Adder_017_io_in2 = io_in[83:78]; // @[RandomHardware.scala 69:41]
  assign Comp_Adder_018_io_in1 = temp_vertex_018[1:0]; // @[RandomHardware.scala 132:51]
  assign Comp_Adder_018_io_in2 = temp_vertex_018[3:2]; // @[RandomHardware.scala 133:51]
  assign Comp_Adder_019_io_in1 = io_in[90:84]; // @[RandomHardware.scala 70:41]
  assign Comp_Adder_019_io_in2 = io_in[97:91]; // @[RandomHardware.scala 71:41]
  assign Comp_Adder_020_io_in1 = temp_vertex_020[3:0]; // @[RandomHardware.scala 98:51]
  assign Comp_Adder_020_io_in2 = temp_vertex_020[7:4]; // @[RandomHardware.scala 99:51]
endmodule
